----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    06:38:45 01/27/2023 
-- Design Name: 
-- Module Name:    halfsubt - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity halfsubt is
    Port ( a : in  STD_LOGIC;
           b : in  STD_LOGIC;
           aa : out  STD_LOGIC;
           bb : out  STD_LOGIC);
end halfsubt;

architecture Behavioral of halfsubt is

begin

process(a,b)

begin
	
	aa <= a xor b;
	
	if(a='0' and b='1')
	then
		bb <= '1';
	else
		bb <= '0';
	end if;

end process;

end Behavioral;

